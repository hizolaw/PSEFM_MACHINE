`ifndef __VECTOR__HEADER__
    `define __VECTOR__HEADER__

    `define RESET_VECTOR    32'hbfc00000
    `define INT_VECTOR    32'hbfc00380
    
`endif
