`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/12/2017 10:48:10 AM
// Design Name: 
// Module Name: time_trigger_tasks
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`include"cp2.vh"
`include"bus.vh"
`include"signal.vh"
module time_trigger_tasks(
    input clk,
    input rst,                  // reset
    input [`TasksNumAddrBus] task_sel,       //要求修改的当前的任务
    input [`TasksNumAddrBus] task_sel_r,       //要求输出的当前的任务
    input [`WORDDATABUS] g_time,//全局时间
    input chs_ena,          //任务状态修改enable
    input new_status,      //新的任务的状态：挂起或就绪
    input [1:0] task_aord_op, //添加/删除任务，高位使能要求操作，低位1为添加，0为删除
    input chcy_ena,   //改变周期掩码使能
    input chph_ena,   //change the phase enable
    input chdeadline_ena,   //change the deadline enable
    input chcyen_ena, //改变是否周期使能
    input cyen_op,
    input [`WORDDATABUS] task_write_data_input,//new phase
    input trigger_op_ena,  //time trigger enable edit enable
    input trigger_op,  // new time tirgger status
    //input [`TasksNumAddrBus] running_task,
//    input time_cy_read_ena,
//    input time_ph_read_ena,
//    input deadline_read_ena,
//    input pri_read_ena,
//    input task_status_read_ena,
//    input task_trigger_read_ena,
    input  [2:0] info_sel,//0:周期信息，1：相位信息，2：死线信息，3：任务是否周期，4：任务时间触发，5：任务状态，6：任务是否存在,7：返回0
    output reg [`WORDADDRBUS] task_info,
    output reg [`TasksNumAddrBusAddOne] tt_top_pri_task,  //top privity task's privity 
    output reg [`TasksNumAddrBusAddOne] et_top_pri_task,  //top privity task's privity 
    //output reg [`TasksNumAddrBusAddOne] second_pri_task,//second privity task's privity 
    output reg [`DoubleWordDataBus] deadline_warn, // when it's high,at least one task arrive deadline
    output wire [`DoubleWordDataBus] task_exist_list_output
    );
    
    reg [`TasksNumAddrBus] deadline_task;
    reg [`DoubleWordDataBus] task_exist_list;
    reg [`DoubleWordDataBus] task_status_list;
    reg [`DoubleWordDataBus] task_cyen_list;
    reg [`DoubleWordDataBus] task_tg_en;
    reg [`DoubleWordDataBus] task_tg_conf;
    reg [`WORDDATABUS] task_tg_cymask[`TR_TASKS_NUM-1:0];
    reg [`WORDDATABUS] task_tg_ph[`TR_TASKS_NUM-1:0];
    reg [`WORDDATABUS] task_tg_deadline[`TR_TASKS_NUM-1:0];
    wire [`DoubleWordDataBus] task_sel_mask;
    assign task_sel_mask = `DOUBLEWORD_DATA_W'b1<<task_sel;
    assign task_exist_list_output=task_exist_list;  
     
    //数据读
    always @(*)begin
        if(rst==`RESET_ENABLE)begin
            task_info=0;
        end else begin
            case (info_sel)
            `PH_INFO:task_info=task_tg_ph[task_sel_r];
            `DEADLINE_INFO:task_info=task_tg_deadline[task_sel_r];
            `STATUS_INFO:task_info=(task_status_list&task_sel_mask)>>task_sel_r;
            `TRIGGER_INFO:task_info=(task_tg_en&task_sel_mask)>>task_sel_r;
            `IS_CY_INFO:task_info=(task_cyen_list&task_sel_mask)>>task_sel_r;
            `CY_INFO:task_info=task_tg_cymask[task_sel_r];
            default:task_info=0;
            endcase
        end
    end
    //deadline的设置
    always @(posedge clk or `RESET_EDGE rst)begin
        if(rst==`RESET_ENABLE)begin
            task_tg_deadline[0]<=`WORD_DATA_W'b0;
            task_tg_deadline[1]<=`WORD_DATA_W'b0;
            task_tg_deadline[2]<=`WORD_DATA_W'b0;
            task_tg_deadline[3]<=`WORD_DATA_W'b0;
            task_tg_deadline[4]<=`WORD_DATA_W'b0;
            task_tg_deadline[5]<=`WORD_DATA_W'b0;
            task_tg_deadline[6]<=`WORD_DATA_W'b0;
            task_tg_deadline[7]<=`WORD_DATA_W'b0;
            task_tg_deadline[8]<=`WORD_DATA_W'b0;
            task_tg_deadline[9]<=`WORD_DATA_W'b0;
            task_tg_deadline[10]<=`WORD_DATA_W'b0;
            task_tg_deadline[11]<=`WORD_DATA_W'b0;
            task_tg_deadline[12]<=`WORD_DATA_W'b0;
            task_tg_deadline[13]<=`WORD_DATA_W'b0;
            task_tg_deadline[14]<=`WORD_DATA_W'b0;
            task_tg_deadline[15]<=`WORD_DATA_W'b0;
            task_tg_deadline[16]<=`WORD_DATA_W'b0;
            task_tg_deadline[17]<=`WORD_DATA_W'b0;
            task_tg_deadline[18]<=`WORD_DATA_W'b0;
            task_tg_deadline[19]<=`WORD_DATA_W'b0;
            task_tg_deadline[20]<=`WORD_DATA_W'b0;
            task_tg_deadline[21]<=`WORD_DATA_W'b0;
            task_tg_deadline[22]<=`WORD_DATA_W'b0;
            task_tg_deadline[23]<=`WORD_DATA_W'b0;
            task_tg_deadline[24]<=`WORD_DATA_W'b0;
            task_tg_deadline[25]<=`WORD_DATA_W'b0;
            task_tg_deadline[26]<=`WORD_DATA_W'b0;
            task_tg_deadline[27]<=`WORD_DATA_W'b0;
            task_tg_deadline[28]<=`WORD_DATA_W'b0;
            task_tg_deadline[29]<=`WORD_DATA_W'b0;
            task_tg_deadline[30]<=`WORD_DATA_W'b0;
            task_tg_deadline[31]<=`WORD_DATA_W'b0;
            task_tg_deadline[32]<=`WORD_DATA_W'b0;
            task_tg_deadline[33]<=`WORD_DATA_W'b0;
            task_tg_deadline[34]<=`WORD_DATA_W'b0;
            task_tg_deadline[35]<=`WORD_DATA_W'b0;
            task_tg_deadline[36]<=`WORD_DATA_W'b0;
            task_tg_deadline[37]<=`WORD_DATA_W'b0;
            task_tg_deadline[38]<=`WORD_DATA_W'b0;
            task_tg_deadline[39]<=`WORD_DATA_W'b0;
            task_tg_deadline[40]<=`WORD_DATA_W'b0;
            task_tg_deadline[41]<=`WORD_DATA_W'b0;
            task_tg_deadline[42]<=`WORD_DATA_W'b0;
            task_tg_deadline[43]<=`WORD_DATA_W'b0;
            task_tg_deadline[44]<=`WORD_DATA_W'b0;
            task_tg_deadline[45]<=`WORD_DATA_W'b0;
            task_tg_deadline[46]<=`WORD_DATA_W'b0;
            task_tg_deadline[47]<=`WORD_DATA_W'b0;
            task_tg_deadline[48]<=`WORD_DATA_W'b0;
            task_tg_deadline[49]<=`WORD_DATA_W'b0;
            task_tg_deadline[50]<=`WORD_DATA_W'b0;
            task_tg_deadline[51]<=`WORD_DATA_W'b0;
            task_tg_deadline[52]<=`WORD_DATA_W'b0;
            task_tg_deadline[53]<=`WORD_DATA_W'b0;
            task_tg_deadline[54]<=`WORD_DATA_W'b0;
            task_tg_deadline[55]<=`WORD_DATA_W'b0;
            task_tg_deadline[56]<=`WORD_DATA_W'b0;
            task_tg_deadline[57]<=`WORD_DATA_W'b0;
            task_tg_deadline[58]<=`WORD_DATA_W'b0;
            task_tg_deadline[59]<=`WORD_DATA_W'b0;
            task_tg_deadline[60]<=`WORD_DATA_W'b0;
            task_tg_deadline[61]<=`WORD_DATA_W'b0;
            task_tg_deadline[62]<=`WORD_DATA_W'b0;
            task_tg_deadline[63]<=`WORD_DATA_W'b0;
        end else begin
            if(chdeadline_ena)begin
                task_tg_deadline[task_sel]<=task_write_data_input+task_tg_ph[task_sel];
            end
        end
    end


    //任务时间触发使能和关闭
    always @(posedge clk or `RESET_EDGE rst)begin
        if(rst==`RESET_ENABLE)begin
            task_tg_en<=0;
        end else begin
            if(trigger_op_ena)begin
                task_tg_en<=(trigger_op)?task_tg_en|task_sel_mask:task_tg_en&(~task_sel_mask);
            end else begin
                task_tg_en<=task_tg_en^(task_status_list&(~task_cyen_list));
            end
        end
    end
    //deadline检查
    always @(posedge clk or `RESET_EDGE rst)begin
        if(rst==`RESET_ENABLE)begin
            deadline_warn<=`DOUBLEWORD_DATA_W'b0;
        end else begin
            deadline_warn[0:0]<=task_exist_list[0:0]?
            	((((g_time&task_tg_cymask[0])==task_tg_deadline[0])&&task_status_list[0:0])?
            		1:
            		0):
            	0;
            deadline_warn[1:1]<=task_exist_list[1:1]?
            	((((g_time&task_tg_cymask[1])==task_tg_deadline[1])&&task_status_list[1:1])?
            		1:
            		0):
            	0;
            deadline_warn[2:2]<=task_exist_list[2:2]?
            	((((g_time&task_tg_cymask[2])==task_tg_deadline[2])&&task_status_list[2:2])?
            		1:
            		0):
            	0;
            deadline_warn[3:3]<=task_exist_list[3:3]?
            	((((g_time&task_tg_cymask[3])==task_tg_deadline[3])&&task_status_list[3:3])?
            		1:
            		0):
            	0;
            deadline_warn[4:4]<=task_exist_list[4:4]?
            	((((g_time&task_tg_cymask[4])==task_tg_deadline[4])&&task_status_list[4:4])?
            		1:
            		0):
            	0;
            deadline_warn[5:5]<=task_exist_list[5:5]?
            	((((g_time&task_tg_cymask[5])==task_tg_deadline[5])&&task_status_list[5:5])?
            		1:
            		0):
            	0;
            deadline_warn[6:6]<=task_exist_list[6:6]?
            	((((g_time&task_tg_cymask[6])==task_tg_deadline[6])&&task_status_list[6:6])?
            		1:
            		0):
            	0;
            deadline_warn[7:7]<=task_exist_list[7:7]?
            	((((g_time&task_tg_cymask[7])==task_tg_deadline[7])&&task_status_list[7:7])?
            		1:
            		0):
            	0;
            deadline_warn[8:8]<=task_exist_list[8:8]?
            	((((g_time&task_tg_cymask[8])==task_tg_deadline[8])&&task_status_list[8:8])?
            		1:
            		0):
            	0;
            deadline_warn[9:9]<=task_exist_list[9:9]?
            	((((g_time&task_tg_cymask[9])==task_tg_deadline[9])&&task_status_list[9:9])?
            		1:
            		0):
            	0;
            deadline_warn[10:10]<=task_exist_list[10:10]?
            	((((g_time&task_tg_cymask[10])==task_tg_deadline[10])&&task_status_list[10:10])?
            		1:
            		0):
            	0;
            deadline_warn[11:11]<=task_exist_list[11:11]?
            	((((g_time&task_tg_cymask[11])==task_tg_deadline[11])&&task_status_list[11:11])?
            		1:
            		0):
            	0;
            deadline_warn[12:12]<=task_exist_list[12:12]?
            	((((g_time&task_tg_cymask[12])==task_tg_deadline[12])&&task_status_list[12:12])?
            		1:
            		0):
            	0;
            deadline_warn[13:13]<=task_exist_list[13:13]?
            	((((g_time&task_tg_cymask[13])==task_tg_deadline[13])&&task_status_list[13:13])?
            		1:
            		0):
            	0;
            deadline_warn[14:14]<=task_exist_list[14:14]?
            	((((g_time&task_tg_cymask[14])==task_tg_deadline[14])&&task_status_list[14:14])?
            		1:
            		0):
            	0;
            deadline_warn[15:15]<=task_exist_list[15:15]?
            	((((g_time&task_tg_cymask[15])==task_tg_deadline[15])&&task_status_list[15:15])?
            		1:
            		0):
            	0;
            deadline_warn[16:16]<=task_exist_list[16:16]?
            	((((g_time&task_tg_cymask[16])==task_tg_deadline[16])&&task_status_list[16:16])?
            		1:
            		0):
            	0;
            deadline_warn[17:17]<=task_exist_list[17:17]?
            	((((g_time&task_tg_cymask[17])==task_tg_deadline[17])&&task_status_list[17:17])?
            		1:
            		0):
            	0;
            deadline_warn[18:18]<=task_exist_list[18:18]?
            	((((g_time&task_tg_cymask[18])==task_tg_deadline[18])&&task_status_list[18:18])?
            		1:
            		0):
            	0;
            deadline_warn[19:19]<=task_exist_list[19:19]?
            	((((g_time&task_tg_cymask[19])==task_tg_deadline[19])&&task_status_list[19:19])?
            		1:
            		0):
            	0;
            deadline_warn[20:20]<=task_exist_list[20:20]?
            	((((g_time&task_tg_cymask[20])==task_tg_deadline[20])&&task_status_list[20:20])?
            		1:
            		0):
            	0;
            deadline_warn[21:21]<=task_exist_list[21:21]?
            	((((g_time&task_tg_cymask[21])==task_tg_deadline[21])&&task_status_list[21:21])?
            		1:
            		0):
            	0;
            deadline_warn[22:22]<=task_exist_list[22:22]?
            	((((g_time&task_tg_cymask[22])==task_tg_deadline[22])&&task_status_list[22:22])?
            		1:
            		0):
            	0;
            deadline_warn[23:23]<=task_exist_list[23:23]?
            	((((g_time&task_tg_cymask[23])==task_tg_deadline[23])&&task_status_list[23:23])?
            		1:
            		0):
            	0;
            deadline_warn[24:24]<=task_exist_list[24:24]?
            	((((g_time&task_tg_cymask[24])==task_tg_deadline[24])&&task_status_list[24:24])?
            		1:
            		0):
            	0;
            deadline_warn[25:25]<=task_exist_list[25:25]?
            	((((g_time&task_tg_cymask[25])==task_tg_deadline[25])&&task_status_list[25:25])?
            		1:
            		0):
            	0;
            deadline_warn[26:26]<=task_exist_list[26:26]?
            	((((g_time&task_tg_cymask[26])==task_tg_deadline[26])&&task_status_list[26:26])?
            		1:
            		0):
            	0;
            deadline_warn[27:27]<=task_exist_list[27:27]?
            	((((g_time&task_tg_cymask[27])==task_tg_deadline[27])&&task_status_list[27:27])?
            		1:
            		0):
            	0;
            deadline_warn[28:28]<=task_exist_list[28:28]?
            	((((g_time&task_tg_cymask[28])==task_tg_deadline[28])&&task_status_list[28:28])?
            		1:
            		0):
            	0;
            deadline_warn[29:29]<=task_exist_list[29:29]?
            	((((g_time&task_tg_cymask[29])==task_tg_deadline[29])&&task_status_list[29:29])?
            		1:
            		0):
            	0;
            deadline_warn[30:30]<=task_exist_list[30:30]?
            	((((g_time&task_tg_cymask[30])==task_tg_deadline[30])&&task_status_list[30:30])?
            		1:
            		0):
            	0;
            deadline_warn[31:31]<=task_exist_list[31:31]?
            	((((g_time&task_tg_cymask[31])==task_tg_deadline[31])&&task_status_list[31:31])?
            		1:
            		0):
            	0;
            deadline_warn[32:32]<=task_exist_list[32:32]?
            	((((g_time&task_tg_cymask[32])==task_tg_deadline[32])&&task_status_list[32:32])?
            		1:
            		0):
            	0;
            deadline_warn[33:33]<=task_exist_list[33:33]?
            	((((g_time&task_tg_cymask[33])==task_tg_deadline[33])&&task_status_list[33:33])?
            		1:
            		0):
            	0;
            deadline_warn[34:34]<=task_exist_list[34:34]?
            	((((g_time&task_tg_cymask[34])==task_tg_deadline[34])&&task_status_list[34:34])?
            		1:
            		0):
            	0;
            deadline_warn[35:35]<=task_exist_list[35:35]?
            	((((g_time&task_tg_cymask[35])==task_tg_deadline[35])&&task_status_list[35:35])?
            		1:
            		0):
            	0;
            deadline_warn[36:36]<=task_exist_list[36:36]?
            	((((g_time&task_tg_cymask[36])==task_tg_deadline[36])&&task_status_list[36:36])?
            		1:
            		0):
            	0;
            deadline_warn[37:37]<=task_exist_list[37:37]?
            	((((g_time&task_tg_cymask[37])==task_tg_deadline[37])&&task_status_list[37:37])?
            		1:
            		0):
            	0;
            deadline_warn[38:38]<=task_exist_list[38:38]?
            	((((g_time&task_tg_cymask[38])==task_tg_deadline[38])&&task_status_list[38:38])?
            		1:
            		0):
            	0;
            deadline_warn[39:39]<=task_exist_list[39:39]?
            	((((g_time&task_tg_cymask[39])==task_tg_deadline[39])&&task_status_list[39:39])?
            		1:
            		0):
            	0;
            deadline_warn[40:40]<=task_exist_list[40:40]?
            	((((g_time&task_tg_cymask[40])==task_tg_deadline[40])&&task_status_list[40:40])?
            		1:
            		0):
            	0;
            deadline_warn[41:41]<=task_exist_list[41:41]?
            	((((g_time&task_tg_cymask[41])==task_tg_deadline[41])&&task_status_list[41:41])?
            		1:
            		0):
            	0;
            deadline_warn[42:42]<=task_exist_list[42:42]?
            	((((g_time&task_tg_cymask[42])==task_tg_deadline[42])&&task_status_list[42:42])?
            		1:
            		0):
            	0;
            deadline_warn[43:43]<=task_exist_list[43:43]?
            	((((g_time&task_tg_cymask[43])==task_tg_deadline[43])&&task_status_list[43:43])?
            		1:
            		0):
            	0;
            deadline_warn[44:44]<=task_exist_list[44:44]?
            	((((g_time&task_tg_cymask[44])==task_tg_deadline[44])&&task_status_list[44:44])?
            		1:
            		0):
            	0;
            deadline_warn[45:45]<=task_exist_list[45:45]?
            	((((g_time&task_tg_cymask[45])==task_tg_deadline[45])&&task_status_list[45:45])?
            		1:
            		0):
            	0;
            deadline_warn[46:46]<=task_exist_list[46:46]?
            	((((g_time&task_tg_cymask[46])==task_tg_deadline[46])&&task_status_list[46:46])?
            		1:
            		0):
            	0;
            deadline_warn[47:47]<=task_exist_list[47:47]?
            	((((g_time&task_tg_cymask[47])==task_tg_deadline[47])&&task_status_list[47:47])?
            		1:
            		0):
            	0;
            deadline_warn[48:48]<=task_exist_list[48:48]?
            	((((g_time&task_tg_cymask[48])==task_tg_deadline[48])&&task_status_list[48:48])?
            		1:
            		0):
            	0;
            deadline_warn[49:49]<=task_exist_list[49:49]?
            	((((g_time&task_tg_cymask[49])==task_tg_deadline[49])&&task_status_list[49:49])?
            		1:
            		0):
            	0;
            deadline_warn[50:50]<=task_exist_list[50:50]?
            	((((g_time&task_tg_cymask[50])==task_tg_deadline[50])&&task_status_list[50:50])?
            		1:
            		0):
            	0;
            deadline_warn[51:51]<=task_exist_list[51:51]?
            	((((g_time&task_tg_cymask[51])==task_tg_deadline[51])&&task_status_list[51:51])?
            		1:
            		0):
            	0;
            deadline_warn[52:52]<=task_exist_list[52:52]?
            	((((g_time&task_tg_cymask[52])==task_tg_deadline[52])&&task_status_list[52:52])?
            		1:
            		0):
            	0;
            deadline_warn[53:53]<=task_exist_list[53:53]?
            	((((g_time&task_tg_cymask[53])==task_tg_deadline[53])&&task_status_list[53:53])?
            		1:
            		0):
            	0;
            deadline_warn[54:54]<=task_exist_list[54:54]?
            	((((g_time&task_tg_cymask[54])==task_tg_deadline[54])&&task_status_list[54:54])?
            		1:
            		0):
            	0;
            deadline_warn[55:55]<=task_exist_list[55:55]?
            	((((g_time&task_tg_cymask[55])==task_tg_deadline[55])&&task_status_list[55:55])?
            		1:
            		0):
            	0;
            deadline_warn[56:56]<=task_exist_list[56:56]?
            	((((g_time&task_tg_cymask[56])==task_tg_deadline[56])&&task_status_list[56:56])?
            		1:
            		0):
            	0;
            deadline_warn[57:57]<=task_exist_list[57:57]?
            	((((g_time&task_tg_cymask[57])==task_tg_deadline[57])&&task_status_list[57:57])?
            		1:
            		0):
            	0;
            deadline_warn[58:58]<=task_exist_list[58:58]?
            	((((g_time&task_tg_cymask[58])==task_tg_deadline[58])&&task_status_list[58:58])?
            		1:
            		0):
            	0;
            deadline_warn[59:59]<=task_exist_list[59:59]?
            	((((g_time&task_tg_cymask[59])==task_tg_deadline[59])&&task_status_list[59:59])?
            		1:
            		0):
            	0;
            deadline_warn[60:60]<=task_exist_list[60:60]?
            	((((g_time&task_tg_cymask[60])==task_tg_deadline[60])&&task_status_list[60:60])?
            		1:
            		0):
            	0;
            deadline_warn[61:61]<=task_exist_list[61:61]?
            	((((g_time&task_tg_cymask[61])==task_tg_deadline[61])&&task_status_list[61:61])?
            		1:
            		0):
            	0;
            deadline_warn[62:62]<=task_exist_list[62:62]?
            	((((g_time&task_tg_cymask[62])==task_tg_deadline[62])&&task_status_list[62:62])?
            		1:
            		0):
            	0;
            deadline_warn[63:63]<=task_exist_list[63:63]?
            	((((g_time&task_tg_cymask[63])==task_tg_deadline[63])&&task_status_list[63:63])?
            		1:
            		0):
            	0;
        end
    end

    //任务周期掩码修改   
    always @(posedge clk or `RESET_EDGE rst)begin
        if(rst==`RESET_ENABLE)begin
            task_tg_cymask[0] <=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[1] <=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[2] <=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[3] <=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[4] <=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[5] <=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[6] <=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[7] <=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[8] <=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[9] <=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[10]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[11]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[12]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[13]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[14]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[15]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[16]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[17]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[18]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[19]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[20]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[21]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[22]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[23]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[24]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[25]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[26]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[27]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[28]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[29]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[30]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[31]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[32]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[33]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[34]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[35]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[36]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[37]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[38]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[39]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[40]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[41]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[42]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[43]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[44]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[45]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[46]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[47]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[48]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[49]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[50]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[51]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[52]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[53]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[54]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[55]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[56]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[57]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[58]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[59]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[60]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[61]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[62]<=`DOUBLEWORD_DATA_W'hffff_ffff;
            task_tg_cymask[63]<=`DOUBLEWORD_DATA_W'hffff_ffff;
        end 
        else begin
            if(chcy_ena)begin
                task_tg_cymask[task_sel]<=(`WORD_DATA_W'b1<<task_write_data_input[5:0])-1;
            end
        end
    end
    
    //任务时间触发的相位赋值
    always @(posedge clk or `RESET_EDGE rst)begin
        if(rst==`RESET_ENABLE)begin
            task_tg_ph[0]<=0;
            task_tg_ph[1]<=0;
            task_tg_ph[2]<=0;
            task_tg_ph[3]<=0;
            task_tg_ph[4]<=0;
            task_tg_ph[5]<=0;
            task_tg_ph[6]<=0;
            task_tg_ph[7]<=0;
            task_tg_ph[8]<=0;
            task_tg_ph[9]<=0;
            task_tg_ph[10]<=0;
            task_tg_ph[11]<=0;
            task_tg_ph[12]<=0;
            task_tg_ph[13]<=0;
            task_tg_ph[14]<=0;
            task_tg_ph[15]<=0;
            task_tg_ph[16]<=0;
            task_tg_ph[17]<=0;
            task_tg_ph[18]<=0;
            task_tg_ph[19]<=0;
            task_tg_ph[20]<=0;
            task_tg_ph[21]<=0;
            task_tg_ph[22]<=0;
            task_tg_ph[23]<=0;
            task_tg_ph[24]<=0;
            task_tg_ph[25]<=0;
            task_tg_ph[26]<=0;
            task_tg_ph[27]<=0;
            task_tg_ph[28]<=0;
            task_tg_ph[29]<=0;
            task_tg_ph[30]<=0;
            task_tg_ph[31]<=0;
            task_tg_ph[32]<=0;
            task_tg_ph[33]<=0;
            task_tg_ph[34]<=0;
            task_tg_ph[35]<=0;
            task_tg_ph[36]<=0;
            task_tg_ph[37]<=0;
            task_tg_ph[38]<=0;
            task_tg_ph[39]<=0;
            task_tg_ph[40]<=0;
            task_tg_ph[41]<=0;
            task_tg_ph[42]<=0;
            task_tg_ph[43]<=0;
            task_tg_ph[44]<=0;
            task_tg_ph[45]<=0;
            task_tg_ph[46]<=0;
            task_tg_ph[47]<=0;
            task_tg_ph[48]<=0;
            task_tg_ph[49]<=0;
            task_tg_ph[50]<=0;
            task_tg_ph[51]<=0;
            task_tg_ph[52]<=0;
            task_tg_ph[53]<=0;
            task_tg_ph[54]<=0;
            task_tg_ph[55]<=0;
            task_tg_ph[56]<=0;
            task_tg_ph[57]<=0;
            task_tg_ph[58]<=0;
            task_tg_ph[59]<=0;
            task_tg_ph[60]<=0;
            task_tg_ph[61]<=0;
            task_tg_ph[62]<=0;
            task_tg_ph[63]<=0;
        end 
        else begin
            if(chph_ena) begin
                task_tg_ph[task_sel]<=task_write_data_input;
            end
        end
    end


    // 添加/删除 任务
    always @(posedge clk or `RESET_EDGE rst)begin
        if(rst==`RESET_ENABLE)begin
            task_exist_list<=`DOUBLEWORD_DATA_W'b0;
        end else begin
            task_exist_list<=(task_aord_op[1:1])?
                (task_aord_op[0:0]?task_exist_list|task_sel_mask:task_exist_list&(~task_sel_mask)):
                task_exist_list;
        end
    end
    
    //是否周期的修改
    always @(posedge clk or `RESET_EDGE rst)begin
        if(rst==`RESET_ENABLE)begin
            task_cyen_list<=`DOUBLEWORD_DATA_W'b0;
        end else begin
            if(chcyen_ena)begin
                task_cyen_list<=cyen_op?(task_sel_mask|task_cyen_list):((~task_sel_mask)&task_cyen_list);
            end
        end
    end

    //非周期的时间触发的任务，当被触发一次之后，时间触发关闭
    //always @(*)begin
    //    if(rst==`RESET_ENABLE)begin
    //        task_tg_en=`DOUBLEWORD_DATA_W'b0;
    //    end else begin
    //        task_tg_en=task_tg_en^(task_status_list&(~task_cyen_list));
    //    end
    //end

    //任务的时间触发管理
    always @(posedge clk or `RESET_EDGE rst)begin
        if(rst==`RESET_ENABLE)begin
            task_status_list<=0;
        end else begin
            task_status_list[0:0]<=task_exist_list[0:0]?
            		((chs_ena&&task_sel==0)?
            			new_status:
            			((task_tg_en[0:0]&&((g_time&task_tg_cymask[0])==task_tg_ph[0]))?
            				1:
            				task_status_list[0:0])):
            		0;
            task_status_list[1:1]<=task_exist_list[1:1]?
            		((chs_ena&&task_sel==1)?
            			new_status:
            			((task_tg_en[1:1]&&((g_time&task_tg_cymask[1])==task_tg_ph[1]))?
            				1:
            				task_status_list[1:1])):
            		0;
            task_status_list[2:2]<=task_exist_list[2:2]?
            		((chs_ena&&task_sel==2)?
            			new_status:
            			((task_tg_en[2:2]&&((g_time&task_tg_cymask[2])==task_tg_ph[2]))?
            				1:
            				task_status_list[2:2])):
            		0;
            task_status_list[3:3]<=task_exist_list[3:3]?
            		((chs_ena&&task_sel==3)?
            			new_status:
            			((task_tg_en[3:3]&&((g_time&task_tg_cymask[3])==task_tg_ph[3]))?
            				1:
            				task_status_list[3:3])):
            		0;
            task_status_list[4:4]<=task_exist_list[4:4]?
            		((chs_ena&&task_sel==4)?
            			new_status:
            			((task_tg_en[4:4]&&((g_time&task_tg_cymask[4])==task_tg_ph[4]))?
            				1:
            				task_status_list[4:4])):
            		0;
            task_status_list[5:5]<=task_exist_list[5:5]?
            		((chs_ena&&task_sel==5)?
            			new_status:
            			((task_tg_en[5:5]&&((g_time&task_tg_cymask[5])==task_tg_ph[5]))?
            				1:
            				task_status_list[5:5])):
            		0;
            task_status_list[6:6]<=task_exist_list[6:6]?
            		((chs_ena&&task_sel==6)?
            			new_status:
            			((task_tg_en[6:6]&&((g_time&task_tg_cymask[6])==task_tg_ph[6]))?
            				1:
            				task_status_list[6:6])):
            		0;
            task_status_list[7:7]<=task_exist_list[7:7]?
            		((chs_ena&&task_sel==7)?
            			new_status:
            			((task_tg_en[7:7]&&((g_time&task_tg_cymask[7])==task_tg_ph[7]))?
            				1:
            				task_status_list[7:7])):
            		0;
            task_status_list[8:8]<=task_exist_list[8:8]?
            		((chs_ena&&task_sel==8)?
            			new_status:
            			((task_tg_en[8:8]&&((g_time&task_tg_cymask[8])==task_tg_ph[8]))?
            				1:
            				task_status_list[8:8])):
            		0;
            task_status_list[9:9]<=task_exist_list[9:9]?
            		((chs_ena&&task_sel==9)?
            			new_status:
            			((task_tg_en[9:9]&&((g_time&task_tg_cymask[9])==task_tg_ph[9]))?
            				1:
            				task_status_list[9:9])):
            		0;
            task_status_list[10:10]<=task_exist_list[10:10]?
            		((chs_ena&&task_sel==10)?
            			new_status:
            			((task_tg_en[10:10]&&((g_time&task_tg_cymask[10])==task_tg_ph[10]))?
            				1:
            				task_status_list[10:10])):
            		0;
            task_status_list[11:11]<=task_exist_list[11:11]?
            		((chs_ena&&task_sel==11)?
            			new_status:
            			((task_tg_en[11:11]&&((g_time&task_tg_cymask[11])==task_tg_ph[11]))?
            				1:
            				task_status_list[11:11])):
            		0;
            task_status_list[12:12]<=task_exist_list[12:12]?
            		((chs_ena&&task_sel==12)?
            			new_status:
            			((task_tg_en[12:12]&&((g_time&task_tg_cymask[12])==task_tg_ph[12]))?
            				1:
            				task_status_list[12:12])):
            		0;
            task_status_list[13:13]<=task_exist_list[13:13]?
            		((chs_ena&&task_sel==13)?
            			new_status:
            			((task_tg_en[13:13]&&((g_time&task_tg_cymask[13])==task_tg_ph[13]))?
            				1:
            				task_status_list[13:13])):
            		0;
            task_status_list[14:14]<=task_exist_list[14:14]?
            		((chs_ena&&task_sel==14)?
            			new_status:
            			((task_tg_en[14:14]&&((g_time&task_tg_cymask[14])==task_tg_ph[14]))?
            				1:
            				task_status_list[14:14])):
            		0;
            task_status_list[15:15]<=task_exist_list[15:15]?
            		((chs_ena&&task_sel==15)?
            			new_status:
            			((task_tg_en[15:15]&&((g_time&task_tg_cymask[15])==task_tg_ph[15]))?
            				1:
            				task_status_list[15:15])):
            		0;
            task_status_list[16:16]<=task_exist_list[16:16]?
            		((chs_ena&&task_sel==16)?
            			new_status:
            			((task_tg_en[16:16]&&((g_time&task_tg_cymask[16])==task_tg_ph[16]))?
            				1:
            				task_status_list[16:16])):
            		0;
            task_status_list[17:17]<=task_exist_list[17:17]?
            		((chs_ena&&task_sel==17)?
            			new_status:
            			((task_tg_en[17:17]&&((g_time&task_tg_cymask[17])==task_tg_ph[17]))?
            				1:
            				task_status_list[17:17])):
            		0;
            task_status_list[18:18]<=task_exist_list[18:18]?
            		((chs_ena&&task_sel==18)?
            			new_status:
            			((task_tg_en[18:18]&&((g_time&task_tg_cymask[18])==task_tg_ph[18]))?
            				1:
            				task_status_list[18:18])):
            		0;
            task_status_list[19:19]<=task_exist_list[19:19]?
            		((chs_ena&&task_sel==19)?
            			new_status:
            			((task_tg_en[19:19]&&((g_time&task_tg_cymask[19])==task_tg_ph[19]))?
            				1:
            				task_status_list[19:19])):
            		0;
            task_status_list[20:20]<=task_exist_list[20:20]?
            		((chs_ena&&task_sel==20)?
            			new_status:
            			((task_tg_en[20:20]&&((g_time&task_tg_cymask[20])==task_tg_ph[20]))?
            				1:
            				task_status_list[20:20])):
            		0;
            task_status_list[21:21]<=task_exist_list[21:21]?
            		((chs_ena&&task_sel==21)?
            			new_status:
            			((task_tg_en[21:21]&&((g_time&task_tg_cymask[21])==task_tg_ph[21]))?
            				1:
            				task_status_list[21:21])):
            		0;
            task_status_list[22:22]<=task_exist_list[22:22]?
            		((chs_ena&&task_sel==22)?
            			new_status:
            			((task_tg_en[22:22]&&((g_time&task_tg_cymask[22])==task_tg_ph[22]))?
            				1:
            				task_status_list[22:22])):
            		0;
            task_status_list[23:23]<=task_exist_list[23:23]?
            		((chs_ena&&task_sel==23)?
            			new_status:
            			((task_tg_en[23:23]&&((g_time&task_tg_cymask[23])==task_tg_ph[23]))?
            				1:
            				task_status_list[23:23])):
            		0;
            task_status_list[24:24]<=task_exist_list[24:24]?
            		((chs_ena&&task_sel==24)?
            			new_status:
            			((task_tg_en[24:24]&&((g_time&task_tg_cymask[24])==task_tg_ph[24]))?
            				1:
            				task_status_list[24:24])):
            		0;
            task_status_list[25:25]<=task_exist_list[25:25]?
            		((chs_ena&&task_sel==25)?
            			new_status:
            			((task_tg_en[25:25]&&((g_time&task_tg_cymask[25])==task_tg_ph[25]))?
            				1:
            				task_status_list[25:25])):
            		0;
            task_status_list[26:26]<=task_exist_list[26:26]?
            		((chs_ena&&task_sel==26)?
            			new_status:
            			((task_tg_en[26:26]&&((g_time&task_tg_cymask[26])==task_tg_ph[26]))?
            				1:
            				task_status_list[26:26])):
            		0;
            task_status_list[27:27]<=task_exist_list[27:27]?
            		((chs_ena&&task_sel==27)?
            			new_status:
            			((task_tg_en[27:27]&&((g_time&task_tg_cymask[27])==task_tg_ph[27]))?
            				1:
            				task_status_list[27:27])):
            		0;
            task_status_list[28:28]<=task_exist_list[28:28]?
            		((chs_ena&&task_sel==28)?
            			new_status:
            			((task_tg_en[28:28]&&((g_time&task_tg_cymask[28])==task_tg_ph[28]))?
            				1:
            				task_status_list[28:28])):
            		0;
            task_status_list[29:29]<=task_exist_list[29:29]?
            		((chs_ena&&task_sel==29)?
            			new_status:
            			((task_tg_en[29:29]&&((g_time&task_tg_cymask[29])==task_tg_ph[29]))?
            				1:
            				task_status_list[29:29])):
            		0;
            task_status_list[30:30]<=task_exist_list[30:30]?
            		((chs_ena&&task_sel==30)?
            			new_status:
            			((task_tg_en[30:30]&&((g_time&task_tg_cymask[30])==task_tg_ph[30]))?
            				1:
            				task_status_list[30:30])):
            		0;
            task_status_list[31:31]<=task_exist_list[31:31]?
            		((chs_ena&&task_sel==31)?
            			new_status:
            			((task_tg_en[31:31]&&((g_time&task_tg_cymask[31])==task_tg_ph[31]))?
            				1:
            				task_status_list[31:31])):
            		0;
            task_status_list[32:32]<=task_exist_list[32:32]?
            		((chs_ena&&task_sel==32)?
            			new_status:
            			((task_tg_en[32:32]&&((g_time&task_tg_cymask[32])==task_tg_ph[32]))?
            				1:
            				task_status_list[32:32])):
            		0;
            task_status_list[33:33]<=task_exist_list[33:33]?
            		((chs_ena&&task_sel==33)?
            			new_status:
            			((task_tg_en[33:33]&&((g_time&task_tg_cymask[33])==task_tg_ph[33]))?
            				1:
            				task_status_list[33:33])):
            		0;
            task_status_list[34:34]<=task_exist_list[34:34]?
            		((chs_ena&&task_sel==34)?
            			new_status:
            			((task_tg_en[34:34]&&((g_time&task_tg_cymask[34])==task_tg_ph[34]))?
            				1:
            				task_status_list[34:34])):
            		0;
            task_status_list[35:35]<=task_exist_list[35:35]?
            		((chs_ena&&task_sel==35)?
            			new_status:
            			((task_tg_en[35:35]&&((g_time&task_tg_cymask[35])==task_tg_ph[35]))?
            				1:
            				task_status_list[35:35])):
            		0;
            task_status_list[36:36]<=task_exist_list[36:36]?
            		((chs_ena&&task_sel==36)?
            			new_status:
            			((task_tg_en[36:36]&&((g_time&task_tg_cymask[36])==task_tg_ph[36]))?
            				1:
            				task_status_list[36:36])):
            		0;
            task_status_list[37:37]<=task_exist_list[37:37]?
            		((chs_ena&&task_sel==37)?
            			new_status:
            			((task_tg_en[37:37]&&((g_time&task_tg_cymask[37])==task_tg_ph[37]))?
            				1:
            				task_status_list[37:37])):
            		0;
            task_status_list[38:38]<=task_exist_list[38:38]?
            		((chs_ena&&task_sel==38)?
            			new_status:
            			((task_tg_en[38:38]&&((g_time&task_tg_cymask[38])==task_tg_ph[38]))?
            				1:
            				task_status_list[38:38])):
            		0;
            task_status_list[39:39]<=task_exist_list[39:39]?
            		((chs_ena&&task_sel==39)?
            			new_status:
            			((task_tg_en[39:39]&&((g_time&task_tg_cymask[39])==task_tg_ph[39]))?
            				1:
            				task_status_list[39:39])):
            		0;
            task_status_list[40:40]<=task_exist_list[40:40]?
            		((chs_ena&&task_sel==40)?
            			new_status:
            			((task_tg_en[40:40]&&((g_time&task_tg_cymask[40])==task_tg_ph[40]))?
            				1:
            				task_status_list[40:40])):
            		0;
            task_status_list[41:41]<=task_exist_list[41:41]?
            		((chs_ena&&task_sel==41)?
            			new_status:
            			((task_tg_en[41:41]&&((g_time&task_tg_cymask[41])==task_tg_ph[41]))?
            				1:
            				task_status_list[41:41])):
            		0;
            task_status_list[42:42]<=task_exist_list[42:42]?
            		((chs_ena&&task_sel==42)?
            			new_status:
            			((task_tg_en[42:42]&&((g_time&task_tg_cymask[42])==task_tg_ph[42]))?
            				1:
            				task_status_list[42:42])):
            		0;
            task_status_list[43:43]<=task_exist_list[43:43]?
            		((chs_ena&&task_sel==43)?
            			new_status:
            			((task_tg_en[43:43]&&((g_time&task_tg_cymask[43])==task_tg_ph[43]))?
            				1:
            				task_status_list[43:43])):
            		0;
            task_status_list[44:44]<=task_exist_list[44:44]?
            		((chs_ena&&task_sel==44)?
            			new_status:
            			((task_tg_en[44:44]&&((g_time&task_tg_cymask[44])==task_tg_ph[44]))?
            				1:
            				task_status_list[44:44])):
            		0;
            task_status_list[45:45]<=task_exist_list[45:45]?
            		((chs_ena&&task_sel==45)?
            			new_status:
            			((task_tg_en[45:45]&&((g_time&task_tg_cymask[45])==task_tg_ph[45]))?
            				1:
            				task_status_list[45:45])):
            		0;
            task_status_list[46:46]<=task_exist_list[46:46]?
            		((chs_ena&&task_sel==46)?
            			new_status:
            			((task_tg_en[46:46]&&((g_time&task_tg_cymask[46])==task_tg_ph[46]))?
            				1:
            				task_status_list[46:46])):
            		0;
            task_status_list[47:47]<=task_exist_list[47:47]?
            		((chs_ena&&task_sel==47)?
            			new_status:
            			((task_tg_en[47:47]&&((g_time&task_tg_cymask[47])==task_tg_ph[47]))?
            				1:
            				task_status_list[47:47])):
            		0;
            task_status_list[48:48]<=task_exist_list[48:48]?
            		((chs_ena&&task_sel==48)?
            			new_status:
            			((task_tg_en[48:48]&&((g_time&task_tg_cymask[48])==task_tg_ph[48]))?
            				1:
            				task_status_list[48:48])):
            		0;
            task_status_list[49:49]<=task_exist_list[49:49]?
            		((chs_ena&&task_sel==49)?
            			new_status:
            			((task_tg_en[49:49]&&((g_time&task_tg_cymask[49])==task_tg_ph[49]))?
            				1:
            				task_status_list[49:49])):
            		0;
            task_status_list[50:50]<=task_exist_list[50:50]?
            		((chs_ena&&task_sel==50)?
            			new_status:
            			((task_tg_en[50:50]&&((g_time&task_tg_cymask[50])==task_tg_ph[50]))?
            				1:
            				task_status_list[50:50])):
            		0;
            task_status_list[51:51]<=task_exist_list[51:51]?
            		((chs_ena&&task_sel==51)?
            			new_status:
            			((task_tg_en[51:51]&&((g_time&task_tg_cymask[51])==task_tg_ph[51]))?
            				1:
            				task_status_list[51:51])):
            		0;
            task_status_list[52:52]<=task_exist_list[52:52]?
            		((chs_ena&&task_sel==52)?
            			new_status:
            			((task_tg_en[52:52]&&((g_time&task_tg_cymask[52])==task_tg_ph[52]))?
            				1:
            				task_status_list[52:52])):
            		0;
            task_status_list[53:53]<=task_exist_list[53:53]?
            		((chs_ena&&task_sel==53)?
            			new_status:
            			((task_tg_en[53:53]&&((g_time&task_tg_cymask[53])==task_tg_ph[53]))?
            				1:
            				task_status_list[53:53])):
            		0;
            task_status_list[54:54]<=task_exist_list[54:54]?
            		((chs_ena&&task_sel==54)?
            			new_status:
            			((task_tg_en[54:54]&&((g_time&task_tg_cymask[54])==task_tg_ph[54]))?
            				1:
            				task_status_list[54:54])):
            		0;
            task_status_list[55:55]<=task_exist_list[55:55]?
            		((chs_ena&&task_sel==55)?
            			new_status:
            			((task_tg_en[55:55]&&((g_time&task_tg_cymask[55])==task_tg_ph[55]))?
            				1:
            				task_status_list[55:55])):
            		0;
            task_status_list[56:56]<=task_exist_list[56:56]?
            		((chs_ena&&task_sel==56)?
            			new_status:
            			((task_tg_en[56:56]&&((g_time&task_tg_cymask[56])==task_tg_ph[56]))?
            				1:
            				task_status_list[56:56])):
            		0;
            task_status_list[57:57]<=task_exist_list[57:57]?
            		((chs_ena&&task_sel==57)?
            			new_status:
            			((task_tg_en[57:57]&&((g_time&task_tg_cymask[57])==task_tg_ph[57]))?
            				1:
            				task_status_list[57:57])):
            		0;
            task_status_list[58:58]<=task_exist_list[58:58]?
            		((chs_ena&&task_sel==58)?
            			new_status:
            			((task_tg_en[58:58]&&((g_time&task_tg_cymask[58])==task_tg_ph[58]))?
            				1:
            				task_status_list[58:58])):
            		0;
            task_status_list[59:59]<=task_exist_list[59:59]?
            		((chs_ena&&task_sel==59)?
            			new_status:
            			((task_tg_en[59:59]&&((g_time&task_tg_cymask[59])==task_tg_ph[59]))?
            				1:
            				task_status_list[59:59])):
            		0;
            task_status_list[60:60]<=task_exist_list[60:60]?
            		((chs_ena&&task_sel==60)?
            			new_status:
            			((task_tg_en[60:60]&&((g_time&task_tg_cymask[60])==task_tg_ph[60]))?
            				1:
            				task_status_list[60:60])):
            		0;
            task_status_list[61:61]<=task_exist_list[61:61]?
            		((chs_ena&&task_sel==61)?
            			new_status:
            			((task_tg_en[61:61]&&((g_time&task_tg_cymask[61])==task_tg_ph[61]))?
            				1:
            				task_status_list[61:61])):
            		0;
            task_status_list[62:62]<=task_exist_list[62:62]?
            		((chs_ena&&task_sel==62)?
            			new_status:
            			((task_tg_en[62:62]&&((g_time&task_tg_cymask[62])==task_tg_ph[62]))?
            				1:
            				task_status_list[62:62])):
            		0;
            task_status_list[63:63]<=task_exist_list[63:63]?
    		        ((chs_ena&&task_sel==63)?
            			new_status:
            			((task_tg_en[63:63]&&((g_time&task_tg_cymask[63])==task_tg_ph[63]))?
            				1:
            				task_status_list[63:63])):
            		0;
        end
    end

    // 时间触发的最高优先级的任务的选择
    always @(*)begin
        if(rst==`RESET_ENABLE)begin
            tt_top_pri_task=64;
        end else begin
            casex(task_status_list&task_tg_en)
                `DOUBLEWORD_DATA_W'b???????????????????????????????????????????????????????????????1:tt_top_pri_task=0;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????????????????????????????????10:tt_top_pri_task=1;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????????????????????????????????100:tt_top_pri_task=2;
                `DOUBLEWORD_DATA_W'b????????????????????????????????????????????????????????????1000:tt_top_pri_task=3;
                `DOUBLEWORD_DATA_W'b???????????????????????????????????????????????????????????10000:tt_top_pri_task=4;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????????????????????????????100000:tt_top_pri_task=5;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????????????????????????????1000000:tt_top_pri_task=6;
                `DOUBLEWORD_DATA_W'b????????????????????????????????????????????????????????10000000:tt_top_pri_task=7;
                `DOUBLEWORD_DATA_W'b???????????????????????????????????????????????????????100000000:tt_top_pri_task=8;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????????????????????????1000000000:tt_top_pri_task=9;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????????????????????????10000000000:tt_top_pri_task=10;
                `DOUBLEWORD_DATA_W'b????????????????????????????????????????????????????100000000000:tt_top_pri_task=11;
                `DOUBLEWORD_DATA_W'b???????????????????????????????????????????????????1000000000000:tt_top_pri_task=12;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????????????????????10000000000000:tt_top_pri_task=13;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????????????????????100000000000000:tt_top_pri_task=14;
                `DOUBLEWORD_DATA_W'b????????????????????????????????????????????????1000000000000000:tt_top_pri_task=15;
                `DOUBLEWORD_DATA_W'b???????????????????????????????????????????????10000000000000000:tt_top_pri_task=16;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????????????????100000000000000000:tt_top_pri_task=17;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????????????????1000000000000000000:tt_top_pri_task=18;
                `DOUBLEWORD_DATA_W'b????????????????????????????????????????????10000000000000000000:tt_top_pri_task=19;
                `DOUBLEWORD_DATA_W'b???????????????????????????????????????????100000000000000000000:tt_top_pri_task=20;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????????????1000000000000000000000:tt_top_pri_task=21;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????????????10000000000000000000000:tt_top_pri_task=22;
                `DOUBLEWORD_DATA_W'b????????????????????????????????????????100000000000000000000000:tt_top_pri_task=23;
                `DOUBLEWORD_DATA_W'b???????????????????????????????????????1000000000000000000000000:tt_top_pri_task=24;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????????10000000000000000000000000:tt_top_pri_task=25;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????????100000000000000000000000000:tt_top_pri_task=26;
                `DOUBLEWORD_DATA_W'b????????????????????????????????????1000000000000000000000000000:tt_top_pri_task=27;
                `DOUBLEWORD_DATA_W'b???????????????????????????????????10000000000000000000000000000:tt_top_pri_task=28;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????100000000000000000000000000000:tt_top_pri_task=29;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????1000000000000000000000000000000:tt_top_pri_task=30;
                `DOUBLEWORD_DATA_W'b????????????????????????????????10000000000000000000000000000000:tt_top_pri_task=31;
                `DOUBLEWORD_DATA_W'b???????????????????????????????100000000000000000000000000000000:tt_top_pri_task=32;
                `DOUBLEWORD_DATA_W'b??????????????????????????????1000000000000000000000000000000000:tt_top_pri_task=33;
                `DOUBLEWORD_DATA_W'b?????????????????????????????10000000000000000000000000000000000:tt_top_pri_task=34;
                `DOUBLEWORD_DATA_W'b????????????????????????????100000000000000000000000000000000000:tt_top_pri_task=35;
                `DOUBLEWORD_DATA_W'b???????????????????????????1000000000000000000000000000000000000:tt_top_pri_task=36;
                `DOUBLEWORD_DATA_W'b??????????????????????????10000000000000000000000000000000000000:tt_top_pri_task=37;
                `DOUBLEWORD_DATA_W'b?????????????????????????100000000000000000000000000000000000000:tt_top_pri_task=38;
                `DOUBLEWORD_DATA_W'b????????????????????????1000000000000000000000000000000000000000:tt_top_pri_task=39;
                `DOUBLEWORD_DATA_W'b???????????????????????10000000000000000000000000000000000000000:tt_top_pri_task=40;
                `DOUBLEWORD_DATA_W'b??????????????????????100000000000000000000000000000000000000000:tt_top_pri_task=41;
                `DOUBLEWORD_DATA_W'b?????????????????????1000000000000000000000000000000000000000000:tt_top_pri_task=42;
                `DOUBLEWORD_DATA_W'b????????????????????10000000000000000000000000000000000000000000:tt_top_pri_task=43;
                `DOUBLEWORD_DATA_W'b???????????????????100000000000000000000000000000000000000000000:tt_top_pri_task=44;
                `DOUBLEWORD_DATA_W'b??????????????????1000000000000000000000000000000000000000000000:tt_top_pri_task=45;
                `DOUBLEWORD_DATA_W'b?????????????????10000000000000000000000000000000000000000000000:tt_top_pri_task=46;
                `DOUBLEWORD_DATA_W'b????????????????100000000000000000000000000000000000000000000000:tt_top_pri_task=47;
                `DOUBLEWORD_DATA_W'b???????????????1000000000000000000000000000000000000000000000000:tt_top_pri_task=48;
                `DOUBLEWORD_DATA_W'b??????????????10000000000000000000000000000000000000000000000000:tt_top_pri_task=49;
                `DOUBLEWORD_DATA_W'b?????????????100000000000000000000000000000000000000000000000000:tt_top_pri_task=50;
                `DOUBLEWORD_DATA_W'b????????????1000000000000000000000000000000000000000000000000000:tt_top_pri_task=51;
                `DOUBLEWORD_DATA_W'b???????????10000000000000000000000000000000000000000000000000000:tt_top_pri_task=52;
                `DOUBLEWORD_DATA_W'b??????????100000000000000000000000000000000000000000000000000000:tt_top_pri_task=53;
                `DOUBLEWORD_DATA_W'b?????????1000000000000000000000000000000000000000000000000000000:tt_top_pri_task=54;
                `DOUBLEWORD_DATA_W'b????????10000000000000000000000000000000000000000000000000000000:tt_top_pri_task=55;
                `DOUBLEWORD_DATA_W'b???????100000000000000000000000000000000000000000000000000000000:tt_top_pri_task=56;
                `DOUBLEWORD_DATA_W'b??????1000000000000000000000000000000000000000000000000000000000:tt_top_pri_task=57;
                `DOUBLEWORD_DATA_W'b?????10000000000000000000000000000000000000000000000000000000000:tt_top_pri_task=58;
                `DOUBLEWORD_DATA_W'b????100000000000000000000000000000000000000000000000000000000000:tt_top_pri_task=59;
                `DOUBLEWORD_DATA_W'b???1000000000000000000000000000000000000000000000000000000000000:tt_top_pri_task=60;
                `DOUBLEWORD_DATA_W'b??10000000000000000000000000000000000000000000000000000000000000:tt_top_pri_task=61;
                `DOUBLEWORD_DATA_W'b?100000000000000000000000000000000000000000000000000000000000000:tt_top_pri_task=62;
                `DOUBLEWORD_DATA_W'b1000000000000000000000000000000000000000000000000000000000000000:tt_top_pri_task=63;            
                default:tt_top_pri_task<=64;
            endcase
        end
    end
    //事件触发的最高优先级的任务
    always @(*)begin
        if(rst==`RESET_ENABLE)begin
            et_top_pri_task=64;
        end else begin
            casex(task_status_list&(~task_tg_en))
                `DOUBLEWORD_DATA_W'b???????????????????????????????????????????????????????????????1:et_top_pri_task=0;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????????????????????????????????10:et_top_pri_task=1;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????????????????????????????????100:et_top_pri_task=2;
                `DOUBLEWORD_DATA_W'b????????????????????????????????????????????????????????????1000:et_top_pri_task=3;
                `DOUBLEWORD_DATA_W'b???????????????????????????????????????????????????????????10000:et_top_pri_task=4;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????????????????????????????100000:et_top_pri_task=5;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????????????????????????????1000000:et_top_pri_task=6;
                `DOUBLEWORD_DATA_W'b????????????????????????????????????????????????????????10000000:et_top_pri_task=7;
                `DOUBLEWORD_DATA_W'b???????????????????????????????????????????????????????100000000:et_top_pri_task=8;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????????????????????????1000000000:et_top_pri_task=9;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????????????????????????10000000000:et_top_pri_task=10;
                `DOUBLEWORD_DATA_W'b????????????????????????????????????????????????????100000000000:et_top_pri_task=11;
                `DOUBLEWORD_DATA_W'b???????????????????????????????????????????????????1000000000000:et_top_pri_task=12;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????????????????????10000000000000:et_top_pri_task=13;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????????????????????100000000000000:et_top_pri_task=14;
                `DOUBLEWORD_DATA_W'b????????????????????????????????????????????????1000000000000000:et_top_pri_task=15;
                `DOUBLEWORD_DATA_W'b???????????????????????????????????????????????10000000000000000:et_top_pri_task=16;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????????????????100000000000000000:et_top_pri_task=17;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????????????????1000000000000000000:et_top_pri_task=18;
                `DOUBLEWORD_DATA_W'b????????????????????????????????????????????10000000000000000000:et_top_pri_task=19;
                `DOUBLEWORD_DATA_W'b???????????????????????????????????????????100000000000000000000:et_top_pri_task=20;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????????????1000000000000000000000:et_top_pri_task=21;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????????????10000000000000000000000:et_top_pri_task=22;
                `DOUBLEWORD_DATA_W'b????????????????????????????????????????100000000000000000000000:et_top_pri_task=23;
                `DOUBLEWORD_DATA_W'b???????????????????????????????????????1000000000000000000000000:et_top_pri_task=24;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????????10000000000000000000000000:et_top_pri_task=25;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????????100000000000000000000000000:et_top_pri_task=26;
                `DOUBLEWORD_DATA_W'b????????????????????????????????????1000000000000000000000000000:et_top_pri_task=27;
                `DOUBLEWORD_DATA_W'b???????????????????????????????????10000000000000000000000000000:et_top_pri_task=28;
                `DOUBLEWORD_DATA_W'b??????????????????????????????????100000000000000000000000000000:et_top_pri_task=29;
                `DOUBLEWORD_DATA_W'b?????????????????????????????????1000000000000000000000000000000:et_top_pri_task=30;
                `DOUBLEWORD_DATA_W'b????????????????????????????????10000000000000000000000000000000:et_top_pri_task=31;
                `DOUBLEWORD_DATA_W'b???????????????????????????????100000000000000000000000000000000:et_top_pri_task=32;
                `DOUBLEWORD_DATA_W'b??????????????????????????????1000000000000000000000000000000000:et_top_pri_task=33;
                `DOUBLEWORD_DATA_W'b?????????????????????????????10000000000000000000000000000000000:et_top_pri_task=34;
                `DOUBLEWORD_DATA_W'b????????????????????????????100000000000000000000000000000000000:et_top_pri_task=35;
                `DOUBLEWORD_DATA_W'b???????????????????????????1000000000000000000000000000000000000:et_top_pri_task=36;
                `DOUBLEWORD_DATA_W'b??????????????????????????10000000000000000000000000000000000000:et_top_pri_task=37;
                `DOUBLEWORD_DATA_W'b?????????????????????????100000000000000000000000000000000000000:et_top_pri_task=38;
                `DOUBLEWORD_DATA_W'b????????????????????????1000000000000000000000000000000000000000:et_top_pri_task=39;
                `DOUBLEWORD_DATA_W'b???????????????????????10000000000000000000000000000000000000000:et_top_pri_task=40;
                `DOUBLEWORD_DATA_W'b??????????????????????100000000000000000000000000000000000000000:et_top_pri_task=41;
                `DOUBLEWORD_DATA_W'b?????????????????????1000000000000000000000000000000000000000000:et_top_pri_task=42;
                `DOUBLEWORD_DATA_W'b????????????????????10000000000000000000000000000000000000000000:et_top_pri_task=43;
                `DOUBLEWORD_DATA_W'b???????????????????100000000000000000000000000000000000000000000:et_top_pri_task=44;
                `DOUBLEWORD_DATA_W'b??????????????????1000000000000000000000000000000000000000000000:et_top_pri_task=45;
                `DOUBLEWORD_DATA_W'b?????????????????10000000000000000000000000000000000000000000000:et_top_pri_task=46;
                `DOUBLEWORD_DATA_W'b????????????????100000000000000000000000000000000000000000000000:et_top_pri_task=47;
                `DOUBLEWORD_DATA_W'b???????????????1000000000000000000000000000000000000000000000000:et_top_pri_task=48;
                `DOUBLEWORD_DATA_W'b??????????????10000000000000000000000000000000000000000000000000:et_top_pri_task=49;
                `DOUBLEWORD_DATA_W'b?????????????100000000000000000000000000000000000000000000000000:et_top_pri_task=50;
                `DOUBLEWORD_DATA_W'b????????????1000000000000000000000000000000000000000000000000000:et_top_pri_task=51;
                `DOUBLEWORD_DATA_W'b???????????10000000000000000000000000000000000000000000000000000:et_top_pri_task=52;
                `DOUBLEWORD_DATA_W'b??????????100000000000000000000000000000000000000000000000000000:et_top_pri_task=53;
                `DOUBLEWORD_DATA_W'b?????????1000000000000000000000000000000000000000000000000000000:et_top_pri_task=54;
                `DOUBLEWORD_DATA_W'b????????10000000000000000000000000000000000000000000000000000000:et_top_pri_task=55;
                `DOUBLEWORD_DATA_W'b???????100000000000000000000000000000000000000000000000000000000:et_top_pri_task=56;
                `DOUBLEWORD_DATA_W'b??????1000000000000000000000000000000000000000000000000000000000:et_top_pri_task=57;
                `DOUBLEWORD_DATA_W'b?????10000000000000000000000000000000000000000000000000000000000:et_top_pri_task=58;
                `DOUBLEWORD_DATA_W'b????100000000000000000000000000000000000000000000000000000000000:et_top_pri_task=59;
                `DOUBLEWORD_DATA_W'b???1000000000000000000000000000000000000000000000000000000000000:et_top_pri_task=60;
                `DOUBLEWORD_DATA_W'b??10000000000000000000000000000000000000000000000000000000000000:et_top_pri_task=61;
                `DOUBLEWORD_DATA_W'b?100000000000000000000000000000000000000000000000000000000000000:et_top_pri_task=62;
                `DOUBLEWORD_DATA_W'b1000000000000000000000000000000000000000000000000000000000000000:et_top_pri_task=63;            
                default:et_top_pri_task<=64;
            endcase
        end
    end

endmodule
