`ifndef __CTRL_HEADER__
    `define __CTRL_HEADER__
    

    `define        CTRL_COUNT     5'd9
    `define        CTRL_COMPARE   5'd11
    `define        CTRL_STATUS    5'd12
    `define        CTRL_COUSE     5'd13
    `define        CTRL_EPC       5'd14
    `define        CTRL_PRID      5'd15

`endif
